-- fpu.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fpu is
	port (
		dataa  : in  std_logic_vector(31 downto 0) := (others => '0'); -- s1.dataa
		datab  : in  std_logic_vector(31 downto 0) := (others => '0'); --   .datab
		n      : in  std_logic_vector(3 downto 0)  := (others => '0'); --   .n
		result : out std_logic_vector(31 downto 0)                     --   .result
	);
end entity fpu;

architecture rtl of fpu is
	component fpoint2_combi is
		generic (
			arithmetic_present : integer := 1;
			comparison_present : integer := 1
		);
		port (
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			n      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- n
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component fpoint2_combi;

begin

	nios_custom_instr_floating_point_2_combi_0 : component fpoint2_combi
		generic map (
			arithmetic_present => 1,
			comparison_present => 1
		)
		port map (
			dataa  => dataa,  -- s1.dataa
			datab  => datab,  --   .datab
			n      => n,      --   .n
			result => result  --   .result
		);

end architecture rtl; -- of fpu

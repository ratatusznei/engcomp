// megafunction wizard: %ALTECC%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altecc_encoder 

// ============================================================
// File Name: l.v
// Megafunction Name(s):
// 			altecc_encoder
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************

//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

module l (
	data,
	q)/* synthesis synthesis_clearbox = 1 */;

	input	[63:0]  data;
	output	[71:0]  q;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX 10"
// Retrieval info: CONSTANT: lpm_pipeline NUMERIC "0"
// Retrieval info: CONSTANT: width_codeword NUMERIC "72"
// Retrieval info: CONSTANT: width_dataword NUMERIC "64"
// Retrieval info: USED_PORT: data 0 0 64 0 INPUT NODEFVAL "data[63..0]"
// Retrieval info: USED_PORT: q 0 0 72 0 OUTPUT NODEFVAL "q[71..0]"
// Retrieval info: CONNECT: @data 0 0 64 0 data 0 0 64 0
// Retrieval info: CONNECT: q 0 0 72 0 @q 0 0 72 0
// Retrieval info: GEN_FILE: TYPE_NORMAL l.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL l.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL l.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL l.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL l_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL l_bb.v TRUE
